library verilog;
use verilog.vl_types.all;
entity spiTB is
end spiTB;
