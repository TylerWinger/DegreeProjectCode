library verilog;
use verilog.vl_types.all;
entity codeWord_MUL_Function is
end codeWord_MUL_Function;
