library verilog;
use verilog.vl_types.all;
entity divideTB is
end divideTB;
