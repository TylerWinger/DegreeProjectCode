library verilog;
use verilog.vl_types.all;
entity HammingEncoding64 is
end HammingEncoding64;
