library verilog;
use verilog.vl_types.all;
entity ck is
end ck;
