library verilog;
use verilog.vl_types.all;
entity RSDecoderOld is
end RSDecoderOld;
