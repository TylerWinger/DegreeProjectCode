library verilog;
use verilog.vl_types.all;
entity encodingDecodingTB is
end encodingDecodingTB;
