library verilog;
use verilog.vl_types.all;
entity encodingTB is
end encodingTB;
