library verilog;
use verilog.vl_types.all;
entity Hamming_TB is
end Hamming_TB;
