library verilog;
use verilog.vl_types.all;
entity writingFileTest is
end writingFileTest;
