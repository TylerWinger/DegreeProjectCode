library verilog;
use verilog.vl_types.all;
entity RSDecoder is
end RSDecoder;
