library verilog;
use verilog.vl_types.all;
entity spi_msg_if_sv_unit is
end spi_msg_if_sv_unit;
