library verilog;
use verilog.vl_types.all;
entity spi_byte_tb is
end spi_byte_tb;
