library verilog;
use verilog.vl_types.all;
entity HammingEncoding_Storage_TB is
end HammingEncoding_Storage_TB;
