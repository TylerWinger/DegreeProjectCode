library verilog;
use verilog.vl_types.all;
entity decodingTB is
end decodingTB;
