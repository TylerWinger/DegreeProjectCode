module Encoding_64TB (
    output reg clk,

);
    
endmodule