
module writingFileTest (
input SW,
output LED
);

assign LED = SW;


initial begin

end
    
endmodule