library verilog;
use verilog.vl_types.all;
entity codeWord is
end codeWord;
