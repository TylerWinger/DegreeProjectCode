library verilog;
use verilog.vl_types.all;
entity noise_test_top_tb is
end noise_test_top_tb;
