library verilog;
use verilog.vl_types.all;
entity HammingDecoding is
end HammingDecoding;
