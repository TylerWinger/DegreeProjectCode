library verilog;
use verilog.vl_types.all;
entity spi_msg_tb is
end spi_msg_tb;
