library verilog;
use verilog.vl_types.all;
entity X_OR is
    port(
        in_1            : in     vl_logic;
        in_2            : in     vl_logic;
        out_1           : out    vl_logic
    );
end X_OR;
