library verilog;
use verilog.vl_types.all;
entity Hamming_64_TB is
end Hamming_64_TB;
