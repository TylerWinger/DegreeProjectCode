library verilog;
use verilog.vl_types.all;
entity codeWordV2 is
end codeWordV2;
