library verilog;
use verilog.vl_types.all;
entity readingFileTest is
end readingFileTest;
